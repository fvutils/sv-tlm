/*
 */
package sv_tlm;
    typedef class tlm_export;
    `include "tlm_port.svh"
    `include "tlm_export.svh"
    `include "tlm_transport_if.svh"

endpackage
