/**
 * tlm_req_rsp_channel.svh
 *
 * Copyright 2024 Matthew Ballance and Contributors
 *
 * Licensed under the Apache License, Version 2.0 (the "License"); you may 
 * not use this file except in compliance with the License.  
 * You may obtain a copy of the License at:
 *
 *   http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software 
 * distributed under the License is distributed on an "AS IS" BASIS, 
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.  
 * See the License for the specific language governing permissions and 
 * limitations under the License.
 *
 * Created on:
 *     Author: 
 */
class tlm_req_rsp_channel #(type REQ, type RSP);

    tlm_export #(tlm_blocking_init_if #(REQ, RSP))      init_export;
    tlm_export #(tlm_blocking_targ_if #(REQ, RSP))      targ_export;

    function new( int req_size=1, int rsp_size=1);
        init_export = new("init_export");
        targ_export = new("targ_export");
    endfunction

endclass

