
module top;
import smoke::*;

initial begin
    test t = new();
    t.run();
end


endmodule