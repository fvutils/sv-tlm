/*
 */
package sv_tlm;
    typedef class tlm_export;
    `include "tlm_port.svh"
    `include "tlm_export.svh"
    `include "tlm_transport_if.svh"
    `include "tlm_blocking_get_if.svh"
    `include "tlm_blocking_put_if.svh"
    `include "tlm_blocking_init_if.svh"
    `include "tlm_blocking_targ_if.svh"

endpackage
